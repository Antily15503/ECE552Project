module cpu(
    input clk, rst_n,
    output [15:0] pc,
    output hlt
);


endmodule