module add_16bit (
    input [15:0] A, B,
    input cin,
    output [3:0] sum,
    output cout
)

endmodule