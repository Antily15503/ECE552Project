module control(
    input [3:0] opcode,
    output [2:0] AluOp,
    output RegDst, Branch, MemRead, MemtoReg, ALUSrc, MemWrite, RegWrite, Jump
);




endmodule