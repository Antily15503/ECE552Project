module ALU (
    input [15:0] ALU_In1, ALU_In2,
    input [3:0] Opcode,
    output [15:0] ALU_Out,
    output Error
);
endmodule;